--recebe como inputs a saida do comparados , o dinheiro e o preço
